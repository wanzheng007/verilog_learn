
`timescale 1ns/1ps

module vlg_design(
	input i_clk,
	input i_rst_n
    );
	

endmodule

