
`timescale 1ns/1ps

module vlg_design(
	input clk,
	input rst_n
    );
	

endmodule

